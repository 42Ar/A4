.SUBCKT RV 1 2 3
R1 1 2 50
R2 2 3 50
.ENDS
