*---------- 2N7002 Spice Model ----------
.SUBCKT N7002 10 20 30 
*     TERMINALS:  D  G  S
M1 1 2 3 3 NMOS L = 1E-006 W = 1E-006 
RD 10 1 0.976 
RS 30 3 0.001 
RG 20 2 160.6 
CGS 2 3 2E-011 
EGD 12 0 2 1 1 
VFB 14 0 0 
FFB 2 1 VFB 1 
CGD 13 14 5.9E-011 
R1 13 0 1 
D1 12 13 DLIM 
DDG 15 14 DCGD 
R2 12 15 1 
D2 15 0 DLIM 
DSD 3 10 DSUB 
.MODEL NMOS NMOS LEVEL = 3 VMAX = 1E+006 ETA = 0 VTO = 2.154 
+ TOX = 6E-008 NSUB = 1E+016 KP = 0.4654 KAPPA = 1E-015 U0 = 400 
.MODEL DCGD D CJO = 1.2E-011 VJ = 0.6 M = 0.6 
.MODEL DSUB D IS = 6.808E-010 N = 1.576 RS = 0.1408 BV = 72 CJO = 8E-012 VJ = 0.8 M = 0.6474 
.MODEL DLIM D IS = 0.0001 
.ENDS
*Diodes N7002 Spice Model v0 Last Revised 2017/2/9