********************************
* Copyright:                   *
* Vishay Intertechnology, Inc. *
********************************
*Jun 23, 2014
*ECN S14-1290, Rev. B
*This document is intended as a SPICE modeling guideline and does not
*constitute a commercial product data sheet.  Designers should refer to the
*appropriate data sheet of the same number for guaranteed specification
*limits.
.SUBCKT Si2300DS D G S 
M1 3 GX S S NMOS W= 434656u L= 0.25u 
M2 S GX S D PMOS W= 434656u L= 2.182e-07 
R1 D 3 3.630e-02 TC=7.226e-03 1.107e-05 
CGS GX S 2.334e-10 
CGD GX D 9.514e-12 
RG G GY 3.2
RTCV 100 S 1e6 TC=1.085e-04 -1.152e-06 
ETCV GX GY 100 200 1 
ITCV S 100 1u 
VTCV 200 S 1 
DBD S D DBD 
**************************************************************** 
.MODEL NMOS NMOS ( LEVEL = 3 TOX = 3e-8 
+ RS = 1.966e-02 KP = 3.368e-05 NSUB = 1.250e+17 
+ KAPPA = 3.810e-02 ETA = 3.202e-04 NFS = 5.144e+11 
+ LD = 0 IS = 0 TPG = 1) 
*************************************************************** 
.MODEL PMOS PMOS ( LEVEL = 3 TOX = 3e-8 
+NSUB = 1.681e+16 IS = 0 TPG = -1 ) 
**************************************************************** 
.MODEL DBD D ( 
+FC = 0.1 TT = 1.301e-08 T_MEASURED = 25 BV = 32 
+RS = 4.112e-02 N = 1.339e+00 IS = 1.749e-09 
+EG = 1.046e+00 XTI = 2.764e-01 TRS1 = 7.466e-04 
+CJO = 1.326e-10 VJ = 4.309e-01 M = 3.495e-01 ) 
.ENDS 
