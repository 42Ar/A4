*SRC=1N5819;DI_1N5819;Diodes;Si;  40.0V  1.00A  3.00us   Diodes Inc. Schottky Barrier Rectifier
.MODEL DI_1N5819 D  ( IS=390n RS=0.115 BV=40.0 IBV=1.00m
+ CJO=203p  M=0.333 N=1.70 TT=4.32u )