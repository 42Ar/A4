***********************************************************
*
* MMBT3904
*
* Nexperia
*
* Switching NPN Transistor
* IC   = 200 mA
* VCEO = 40 V 
* hFE  = 100 - 300 @ 1V/10mA
*
*
*
*
* Package pinning does not match Spice model pinning.
* Package: SOT 23
* 
* Package Pin 1: Base
* Package Pin 2: Emitter
* Package Pin 3: Collector
*
*
* Extraction date (week/year): 25/2014
* Spicemodel includes temperature dependency
*
**********************************************************
*#
.SUBCKT MMBT3904 1 2 3
Q1 1 2 3 MAIN
D1 2 1 DIODE
*
* Diode D1 is dedicated to improve modeling in reverse
* mode of operation and does not reflect a physical device.
* 
.MODEL MAIN NPN
+ IS = 2.612E-015
+ NF = 1.005
+ ISE = 2.958E-015
+ NE = 1.533
+ BF = 169
+ IKF = 0.08351
+ VAF = 53.92
+ NR = 0.9982
+ ISC = 3.177E-016
+ NC = 1.094
+ BR = 2.107
+ IKR = 0.5
+ VAR = 100
+ RB = 114
+ IRB = 0.001
+ RBM = 6.2
+ RE = 0.04181
+ RC = 0.9576
+ XTB = 1.522
+ EG = 1.11
+ XTI = 4.633
+ CJE = 1.032E-011
+ VJE = 0.6333
+ MJE = 0.2056
+ TF = 3.55E-010
+ XTF = 10
+ VTF = 2
+ ITF = 0.3
+ PTF = 0
+ CJC = 3.181E-012
+ VJC = 0.8831
+ MJC = 0.3242
+ XCJC = 1
+ TR = 1.45E-007
+ CJS = 0
+ VJS = 0.75
+ MJS = 0.333
+ FC = 0.78
.MODEL DIODE D
+ IS = 1.82E-013
+ N = 1.042
+ BV = 1000
+ IBV = 0.001
+ RS = 380.9
+ CJO = 0
+ VJ = 1
+ M = 0.5
+ FC = 0
+ TT = 0
+ EG = 1.11
+ XTI = 3
.ENDS
*
