***********************************************************
*
* BC856B
*
* Nexperia
*
* General purpose PNP Transistor
* IC   = 100 mA
* VCEO = 65 V 
* hFE  = 125 - 250 @ 5V/2mA
* 
*
*
*
* Package pinning does not match Spice model pinning.
* Package: SOT 23
* 
* Package Pin 1: Base
* Package Pin 2: Emitter
* Package Pin 3: Collector
* 
*
* Extraction date (week/year): 19/2020
* Spice model includes temperature dependency
*
**********************************************************
*#
* Transistor Q2, Resistor RQ and Diode D are dedicated to improve modeling in quasi
* saturation area and reverse area of operation. They do not reflect physical devices.
*
.SUBCKT BC856B 1 2 3
Q1 1 2 3 MAIN 0.9607
Q2 11 2 3 MAIN 0.03929
RQ 1 11 561.1
D1 1 2 DIODE
*
.MODEL MAIN PNP
+ IS = 1.95E-014
+ NF = 1.022
+ ISE = 1.253E-014
+ NE = 1.577
+ BF = 297.2
+ IKF = 0.0831
+ VAF = 41.13
+ NR = 1.021
+ ISC = 1.791E-016
+ NC = 1.183
+ BR = 10.02
+ IKR = 0.02503
+ VAR = 16.61
+ RB = 220
+ IRB = 2.5E-005
+ RBM = 0.9
+ RE = 1.045
+ RC = 0.2657
+ XTB = 1.28
+ EG = 1.11
+ XTI = 2.944
+ CJE = 1.095E-011
+ VJE = 0.6608
+ MJE = 0.375
+ TF = 1.2E-009
+ XTF = 3
+ VTF = 3.813
+ ITF = 0.1208
+ PTF = 0
+ CJC = 5.88E-012
+ VJC = 0.5428
+ MJC = 0.39
+ XCJC = 0.459
+ TR = 8.8E-008
+ CJS = 0
+ VJS = 0.75
+ MJS = 0.333
+ FC = 0.9501
.MODEL DIODE D
+ IS = 7.703E-015
+ N = 1.146
+ BV = 1000
+ IBV = 0.001
+ RS = 2.826E+004
+ CJO = 0
+ VJ = 1
+ M = 0.5
+ FC = 0
+ TT = 0
+ EG = 1.11
+ XTI = 3
.ENDS
*
